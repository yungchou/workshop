version https://git-lfs.github.com/spec/v1
oid sha256:538562d49b6bd13a245c83c6ae1fd83cb0bcc9bb3877d1d88ca5792d3d91f989
size 258461696
